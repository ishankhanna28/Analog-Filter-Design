* C:\Users\Ishan's PC\Desktop\Sem 4\Projects\LIC\Innovative Project\BandReject\BRF.sch

* Schematics Version 9.2
* Sat Apr 03 21:28:22 2021



** Analysis setup **
.ac DEC 100 30 3k


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "BRF.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
